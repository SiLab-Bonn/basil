/**
 * ------------------------------------------------------------
 * Copyright (c) All rights reserved
 * SiLab, Institute of Physics, University of Bonn
 * ------------------------------------------------------------
 */

`timescale 1ps / 1ps
`default_nettype none

module test_eth(
    input wire RESET_N,
    input wire clkin,

    output wire [3:0] rgmii_txd,
    output wire rgmii_tx_ctl,
    output wire rgmii_txc,
    input wire [3:0] rgmii_rxd,
    input wire rgmii_rx_ctl,
    input wire rgmii_rxc,
    output wire mdio_phy_mdc,
    inout wire mdio_phy_mdio,
    output wire phy_rst_n,

    output wire [7:0] LED
);

localparam VERSION = 8'd0;

wire RST;
wire CLK125_PLL, CLK125_90_PLL;
wire PLL_FEEDBACK, LOCKED;
PLLE2_BASE #(
    .BANDWIDTH("OPTIMIZED"),  // OPTIMIZED, HIGH, LOW
    .CLKFBOUT_MULT(10),       // Multiply value for all CLKOUT, (2-64)
    .CLKFBOUT_PHASE(0.0),     // Phase offset in degrees of CLKFB, (-360.000-360.000).
    .CLKIN1_PERIOD(10.000),      // Input clock period in ns to ps resolution (i.e. 33.333 is 30 MHz).

    .CLKOUT0_DIVIDE(8),     // Divide amount for CLKOUT0 (1-128)
    .CLKOUT0_DUTY_CYCLE(0.5), // Duty cycle for CLKOUT0 (0.001-0.999).
    .CLKOUT0_PHASE(0.0),      // Phase offset for CLKOUT0 (-360.000-360.000).

    .CLKOUT1_DIVIDE(8),     // Divide amount for CLKOUT0 (1-128)
    .CLKOUT1_DUTY_CYCLE(0.5), // Duty cycle for CLKOUT0 (0.001-0.999).
    .CLKOUT1_PHASE(90.0),      // Phase offset for CLKOUT0 (-360.000-360.000).

    .DIVCLK_DIVIDE(1),        // Master division value, (1-56)
    .REF_JITTER1(0.0),        // Reference input jitter in UI, (0.000-0.999).
    .STARTUP_WAIT("FALSE")     // Delay DONE until PLL Locks, ("TRUE"/"FALSE")
) PLLE2_BASE_inst (
    .CLKOUT0(CLK125_PLL),
    .CLKOUT1(CLK125_90_PLL),
    .CLKOUT2(),
    .CLKOUT3(),
    .CLKOUT4(),
    .CLKOUT5(),

    .CLKFBOUT(PLL_FEEDBACK),
    .LOCKED(LOCKED),     // 1-bit output: LOCK

    // Input 100 MHz clock
    .CLKIN1(clkin),

    // Control Ports
    .PWRDWN(0),
    .RST(!RESET_N),

    // Feedback
    .CLKFBIN(PLL_FEEDBACK)
);

wire PLL_FEEDBACK2, LOCKED2;
wire BUS_CLK_PLL;
PLLE2_BASE #(
    .BANDWIDTH("OPTIMIZED"),
    .CLKFBOUT_MULT(16),
    .CLKFBOUT_PHASE(0.0),
    .CLKIN1_PERIOD(10.000),

    .CLKOUT0_DIVIDE(12),
    .CLKOUT0_DUTY_CYCLE(0.5),
    .CLKOUT0_PHASE(0.0),

    .DIVCLK_DIVIDE(1),
    .REF_JITTER1(0.0),
    .STARTUP_WAIT("FALSE")
) PLLE2_BASE_inst_2 (
    .CLKOUT0(BUS_CLK_PLL),
    .CLKOUT1(),
    .CLKOUT2(),
    .CLKOUT3(),
    .CLKOUT4(),
    .CLKOUT5(),

    .CLKFBOUT(PLL_FEEDBACK2),
    .LOCKED(LOCKED2), // 1-bit output: LOCK

    .CLKIN1(clkin),

    .PWRDWN(0),
    .RST(!RESET_N),

    .CLKFBIN(PLL_FEEDBACK2)
);

wire BUS_CLK;
BUFG BUFG_inst_BUS_CLK (.O(BUS_CLK), .I(BUS_CLK_PLL));  // 133.3MHz

assign RST = !RESET_N | !LOCKED | !LOCKED2;


wire gmii_tx_clk;
wire gmii_tx_en;
wire [7:0] gmii_txd;
wire gmii_tx_er;
wire gmii_crs;
wire gmii_col;
wire gmii_rx_clk;
wire gmii_rx_dv;
wire [7:0] gmii_rxd;
wire gmii_rx_er;
wire mdio_gem_mdc;
wire mdio_gem_i;
wire mdio_gem_o;
wire mdio_gem_t;
wire link_status;
wire [1:0] clock_speed;
wire duplex_status;
reg GMII_1000M;

wire MII_TX_CLK, MII_TX_CLK_90;
BUFGMUX GMIIMUX (.O(MII_TX_CLK), .I0(rgmii_rxc), .I1(CLK125_PLL), .S(GMII_1000M));
BUFGMUX GMIIMUX90 (.O(MII_TX_CLK_90), .I0(rgmii_rxc), .I1(CLK125_90_PLL), .S(GMII_1000M));

rgmii_io rgmii (
    .rgmii_txd(rgmii_txd),
    .rgmii_tx_ctl(rgmii_tx_ctl),
    .rgmii_txc(rgmii_txc),

    .rgmii_rxd(rgmii_rxd),
    .rgmii_rx_ctl(rgmii_rx_ctl),

    .gmii_txd_int(gmii_txd),      // Internal gmii_txd signal.
    .gmii_tx_en_int(gmii_tx_en),
    .gmii_tx_er_int(gmii_tx_er),
    .gmii_col_int(gmii_col),
    .gmii_crs_int(gmii_crs),
    .gmii_rxd_reg(gmii_rxd),   // RGMII double data rate data valid.
    .gmii_rx_dv_reg(gmii_rx_dv), // gmii_rx_dv_ibuf registered in IOBs.
    .gmii_rx_er_reg(gmii_rx_er), // gmii_rx_er_ibuf registered in IOBs.

    .eth_link_status(link_status),
    .eth_clock_speed(clock_speed),
    .eth_duplex_status(duplex_status),

                              // FOllowing are generated by DCMs
    .tx_rgmii_clk_int(MII_TX_CLK),     // Internal RGMII transmitter clock.
    .tx_rgmii_clk90_int(MII_TX_CLK_90),   // Internal RGMII transmitter clock w/ 90 deg phase
    .rx_rgmii_clk_int(rgmii_rxc),     // Internal RGMII receiver clock

    .reset(!phy_rst_n)
);

//assign GMII_1000M = &clock_speed;
always@(posedge BUS_CLK or posedge RST)begin
    if (RST) begin
        GMII_1000M <= 1'b0;
    end else begin
        GMII_1000M <= clock_speed[1];
    end
end

// Instantiate tri-state buffer for MDIO
IOBUF i_iobuf_mdio (
    .O(mdio_gem_i),
    .IO(mdio_phy_mdio),
    .I(mdio_gem_o),
    .T(mdio_gem_t)
);

wire EEPROM_CS, EEPROM_SK, EEPROM_DI;
wire TCP_CLOSE_REQ;
wire RBCP_ACT, RBCP_WE, RBCP_RE;
wire [7:0] RBCP_WD, RBCP_RD;
wire [31:0] RBCP_ADDR;
wire TCP_RX_WR;
wire [7:0] TCP_RX_DATA;
//reg  [15:0] TCP_RX_WC;
wire [15:0] TCP_RX_WC;
wire RBCP_ACK;
wire SiTCP_RST;

wire TCP_TX_FULL;
wire TCP_TX_WR;
wire [7:0] TCP_TX_DATA;

WRAP_SiTCP_GMII_XC7K_32K #(
    .TIM_PERIOD(8'd133)
) sitcp (
    .CLK(BUS_CLK)                    ,    // in    : System Clock >129MHz
    .RST(RST)                    ,    // in    : System reset
    // Configuration parameters
    .FORCE_DEFAULTn(1'b0)        ,    // in    : Load default parameters
    .EXT_IP_ADDR(32'hc0a80a10)            ,    // in    : IP address[31:0] //192.168.10.16
    .EXT_TCP_PORT(16'd24)        ,    // in    : TCP port #[15:0]
    .EXT_RBCP_PORT(16'd4660)        ,    // in    : RBCP port #[15:0]
    .PHY_ADDR(5'd3)            ,    // in    : PHY-device MIF address[4:0]
    // EEPROM
    .EEPROM_CS(EEPROM_CS)            ,    // out    : Chip select
    .EEPROM_SK(EEPROM_SK)            ,    // out    : Serial data clock
    .EEPROM_DI(EEPROM_DI)            ,    // out    : Serial write data
    .EEPROM_DO(1'b0)            ,    // in    : Serial read data
    // user data, intialial values are stored in the EEPROM, 0xFFFF_FC3C-3F
    .USR_REG_X3C()            ,    // out    : Stored at 0xFFFF_FF3C
    .USR_REG_X3D()            ,    // out    : Stored at 0xFFFF_FF3D
    .USR_REG_X3E()            ,    // out    : Stored at 0xFFFF_FF3E
    .USR_REG_X3F()            ,    // out    : Stored at 0xFFFF_FF3F
    // MII interface
    .GMII_RSTn(phy_rst_n)            ,    // out    : PHY reset
    .GMII_1000M(GMII_1000M)            ,    // in    : GMII mode (0:MII, 1:GMII)
    // TX
    .GMII_TX_CLK(MII_TX_CLK)            ,    // in    : Tx clock
    .GMII_TX_EN(gmii_tx_en)            ,    // out    : Tx enable
    .GMII_TXD(gmii_txd)            ,    // out    : Tx data[7:0]
    .GMII_TX_ER(gmii_tx_er)            ,    // out    : TX error
    // RX
    .GMII_RX_CLK(rgmii_rxc)           ,    // in    : Rx clock
    .GMII_RX_DV(gmii_rx_dv)            ,    // in    : Rx data valid
    .GMII_RXD(gmii_rxd)            ,    // in    : Rx data[7:0]
    .GMII_RX_ER(gmii_rx_er)            ,    // in    : Rx error
    .GMII_CRS(gmii_crs)            ,    // in    : Carrier sense
    .GMII_COL(gmii_col)            ,    // in    : Collision detected
    // Management IF
    .GMII_MDC(mdio_phy_mdc)            ,    // out    : Clock for MDIO
    .GMII_MDIO_IN(mdio_gem_i)        ,    // in    : Data
    .GMII_MDIO_OUT(mdio_gem_o)        ,    // out    : Data
    .GMII_MDIO_OE(mdio_gem_t)        ,    // out    : MDIO output enable
    // User I/F
    .SiTCP_RST(SiTCP_RST)            ,    // out    : Reset for SiTCP and related circuits
    // TCP connection control
    .TCP_OPEN_REQ(1'b0)        ,    // in    : Reserved input, shoud be 0
    .TCP_OPEN_ACK()        ,    // out    : Acknowledge for open (=Socket busy)
    .TCP_ERROR()            ,    // out    : TCP error, its active period is equal to MSL
    .TCP_CLOSE_REQ(TCP_CLOSE_REQ)        ,    // out    : Connection close request
    .TCP_CLOSE_ACK(TCP_CLOSE_REQ)        ,    // in    : Acknowledge for closing
    // FIFO I/F
    .TCP_RX_WC(TCP_RX_WC)            ,    // in    : Rx FIFO write count[15:0] (Unused bits should be set 1)
    .TCP_RX_WR(TCP_RX_WR)            ,    // out    : Write enable
    .TCP_RX_DATA(TCP_RX_DATA)            ,    // out    : Write data[7:0]
    .TCP_TX_FULL(TCP_TX_FULL)            ,    // out    : Almost full flag
    .TCP_TX_WR(TCP_TX_WR)            ,    // in    : Write enable
    .TCP_TX_DATA(TCP_TX_DATA)            ,    // in    : Write data[7:0]
    // RBCP
    .RBCP_ACT(RBCP_ACT)            ,    // out    : RBCP active
    .RBCP_ADDR(RBCP_ADDR)            ,    // out    : Address[31:0]
    .RBCP_WD(RBCP_WD)                ,    // out    : Data[7:0]
    .RBCP_WE(RBCP_WE)                ,    // out    : Write enable
    .RBCP_RE(RBCP_RE)                ,    // out    : Read enable
    .RBCP_ACK(RBCP_ACK)            ,    // in    : Access acknowledge
    .RBCP_RD(RBCP_RD)                    // in    : Read data[7:0]
);

// -------  BUS SYGNALING  ------- //

wire BUS_WR, BUS_RD, BUS_RST;
wire [31:0] BUS_ADD;
wire [7:0] BUS_DATA;
wire INVALID;
assign BUS_RST = SiTCP_RST;

tcp_to_bus itcp_to_bus (
    .BUS_RST(BUS_RST),
    .BUS_CLK(BUS_CLK),

    .TCP_RX_WC(TCP_RX_WC),
    .TCP_RX_WR(TCP_RX_WR),
    .TCP_RX_DATA(TCP_RX_DATA),

    .RBCP_ACT(RBCP_ACT),
    .RBCP_ADDR(RBCP_ADDR),
    .RBCP_WD(RBCP_WD),
    .RBCP_WE(RBCP_WE),
    .RBCP_RE(RBCP_RE),
    .RBCP_ACK(RBCP_ACK),
    .RBCP_RD(RBCP_RD),

    .BUS_WR(BUS_WR),
    .BUS_RD(BUS_RD),
    .BUS_ADD(BUS_ADD),
    .BUS_DATA(BUS_DATA),

    .INVALID(INVALID)
);

// -------  MODULE ADREESSES  ------- //

// Registers
wire SOFT_RST; // Address: 0
assign SOFT_RST = (BUS_ADD == 0 && BUS_WR);

// reset sync
// when writing to addr = 0 then reset
reg RST_FF, RST_FF2, BUS_RST_FF, BUS_RST_FF2;
always @(posedge BUS_CLK) begin
    RST_FF <= SOFT_RST;
    RST_FF2 <= RST_FF;
    BUS_RST_FF <= BUS_RST;
    BUS_RST_FF2 <= BUS_RST_FF;
end

wire SOFT_RST_FLAG;
assign SOFT_RST_FLAG = ~RST_FF2 & RST_FF;
wire BUS_RST_FLAG;
assign BUS_RST_FLAG = BUS_RST_FF2 & ~BUS_RST_FF; // trailing edge
wire RESET;
assign RESET = BUS_RST_FLAG | SOFT_RST_FLAG;

reg [7:0] status_regs[39:0];

wire [7:0] SETUP;
assign SETUP = status_regs[1];
wire [63:0] TEST_DATA;
assign TEST_DATA = {status_regs[9], status_regs[8], status_regs[7], status_regs[6],status_regs[5], status_regs[4], status_regs[3], status_regs[2]};
wire [15:0] TCP_WRITE_DLY;
assign TCP_WRITE_DLY = {status_regs[15], status_regs[14]};

always @(posedge BUS_CLK)
begin
    if(RESET)
    begin
        status_regs[0] <= 8'b0; // Version, Reset
        status_regs[1] <= 8'b0; // Setup
        status_regs[2] <= 8'b0; // Test data
        status_regs[3] <= 8'b0; // Test data
        status_regs[4] <= 8'b0; // Test data
        status_regs[5] <= 8'b0; // Test data
        status_regs[6] <= 8'b0; // Test data
        status_regs[7] <= 8'b0; // Test data
        status_regs[8] <= 8'b0; // Test data
        status_regs[9] <= 8'b0; // Test data
        status_regs[10] <= 8'b0; // UDP write counter
        status_regs[11] <= 8'b0; // UDP write counter
        status_regs[12] <= 8'b0; // UDP write counter
        status_regs[13] <= 8'b0; // UDP write counter
        status_regs[14] <= 8'b0; // TCP write delay
        status_regs[15] <= 8'b0; // TCP write delay
        status_regs[16] <= 8'b0; // TCP write counter
        status_regs[17] <= 8'b0; // TCP write counter
        status_regs[18] <= 8'b0; // TCP write counter
        status_regs[19] <= 8'b0; // TCP write counter
        status_regs[20] <= 8'b0; // TCP write counter
        status_regs[21] <= 8'b0; // TCP write counter
        status_regs[22] <= 8'b0; // TCP write counter
        status_regs[23] <= 8'b0; // TCP write counter
        status_regs[24] <= 8'b0; // TCP failed write counter
        status_regs[25] <= 8'b0; // TCP failed write counter
        status_regs[26] <= 8'b0; // TCP failed write counter
        status_regs[27] <= 8'b0; // TCP failed write counter
        status_regs[28] <= 8'b0; // TCP failed write counter
        status_regs[29] <= 8'b0; // TCP failed write counter
        status_regs[30] <= 8'b0; // TCP failed write counter
        status_regs[31] <= 8'b0; // TCP failed write counter
        status_regs[32] <= 8'b0; // TCP recv write counter
        status_regs[33] <= 8'b0; // TCP recv write counter
        status_regs[34] <= 8'b0; // TCP recv write counter
        status_regs[35] <= 8'b0; // TCP recv write counter
        status_regs[36] <= 8'b0; // TCP recv write counter
        status_regs[37] <= 8'b0; // TCP recv write counter
        status_regs[38] <= 8'b0; // TCP recv write counter
        status_regs[39] <= 8'b0; // TCP recv write counter
    end
    else if(BUS_WR && BUS_ADD < 40)
    begin
        status_regs[BUS_ADD[5:0]] <= BUS_DATA;
    end
end

reg [31:0] UDP_WRITE_CNT;
reg [63:0] TCP_WRITE_CNT;
reg [63:0] TCP_FAILED_WRITE_CNT;
reg [63:0] TCP_RCV_WRITE_CNT;

reg [7:0] BUS_DATA_OUT;
always @ (posedge BUS_CLK) begin
    if(BUS_RD) begin
        if (BUS_ADD == 0)
            BUS_DATA_OUT <= VERSION[7:0];
        else if (BUS_ADD == 1)
            BUS_DATA_OUT <= SETUP;
        else if (BUS_ADD == 2)
            BUS_DATA_OUT <= TEST_DATA[7:0];
        else if (BUS_ADD == 3)
            BUS_DATA_OUT <= TEST_DATA[15:8];
        else if (BUS_ADD == 4)
            BUS_DATA_OUT <= TEST_DATA[23:16];
        else if (BUS_ADD == 5)
            BUS_DATA_OUT <= TEST_DATA[31:24];
        else if (BUS_ADD == 6)
            BUS_DATA_OUT <= TEST_DATA[39:32];
        else if (BUS_ADD == 7)
            BUS_DATA_OUT <= TEST_DATA[47:40];
        else if (BUS_ADD == 8)
            BUS_DATA_OUT <= TEST_DATA[55:48];
        else if (BUS_ADD == 9)
            BUS_DATA_OUT <= TEST_DATA[63:56];
        else if (BUS_ADD == 10)
            BUS_DATA_OUT <= UDP_WRITE_CNT[7:0];
        else if (BUS_ADD == 11)
            BUS_DATA_OUT <= UDP_WRITE_CNT[15:8];
        else if (BUS_ADD == 12)
            BUS_DATA_OUT <= UDP_WRITE_CNT[23:16];
        else if (BUS_ADD == 13)
            BUS_DATA_OUT <= UDP_WRITE_CNT[31:24];
        else if (BUS_ADD == 14)
            BUS_DATA_OUT <= TCP_WRITE_DLY[7:0];
        else if (BUS_ADD == 15)
            BUS_DATA_OUT <= TCP_WRITE_DLY[15:8];
        else if (BUS_ADD == 16)
            BUS_DATA_OUT <= TCP_WRITE_CNT[7:0];
        else if (BUS_ADD == 17)
            BUS_DATA_OUT <= TCP_WRITE_CNT[15:8];
        else if (BUS_ADD == 18)
            BUS_DATA_OUT <= TCP_WRITE_CNT[23:16];
        else if (BUS_ADD == 19)
            BUS_DATA_OUT <= TCP_WRITE_CNT[31:24];
        else if (BUS_ADD == 20)
            BUS_DATA_OUT <= TCP_WRITE_CNT[39:32];
        else if (BUS_ADD == 21)
            BUS_DATA_OUT <= TCP_WRITE_CNT[47:40];
        else if (BUS_ADD == 22)
            BUS_DATA_OUT <= TCP_WRITE_CNT[55:48];
        else if (BUS_ADD == 23)
            BUS_DATA_OUT <= TCP_WRITE_CNT[63:56];
        else if (BUS_ADD == 24)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[7:0];
        else if (BUS_ADD == 25)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[15:8];
        else if (BUS_ADD == 26)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[23:16];
        else if (BUS_ADD == 27)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[31:24];
        else if (BUS_ADD == 28)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[39:32];
        else if (BUS_ADD == 29)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[47:40];
        else if (BUS_ADD == 30)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[55:48];
        else if (BUS_ADD == 31)
            BUS_DATA_OUT <= TCP_FAILED_WRITE_CNT[63:56];
        else if (BUS_ADD == 32)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[7:0];
        else if (BUS_ADD == 33)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[15:8];
        else if (BUS_ADD == 34)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[23:16];
        else if (BUS_ADD == 35)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[31:24];
        else if (BUS_ADD == 36)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[39:32];
        else if (BUS_ADD == 37)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[47:40];
        else if (BUS_ADD == 38)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[55:48];
        else if (BUS_ADD == 39)
            BUS_DATA_OUT <= TCP_RCV_WRITE_CNT[63:56];
        else
            BUS_DATA_OUT <= 0;
    end
end


reg BUS_READ;
always @ (posedge BUS_CLK)
    if (BUS_RD & BUS_ADD < 40)
        BUS_READ <= 1;
    else
        BUS_READ <= 0;

assign BUS_DATA = BUS_READ ? BUS_DATA_OUT : 8'hzz;

// Test registers

wire recv_tcp_data_wfull;
wire RECV_TCP_DATA_FULL;
assign RECV_TCP_DATA_FULL = recv_tcp_data_wfull;
wire recv_tcp_data_cdc_fifo_write;
assign recv_tcp_data_cdc_fifo_write = 1'b0; //TCP_RX_WR & ~RECV_TCP_DATA_FULL;
wire recv_tcp_data_fifo_full, recv_tcp_data_cdc_fifo_empty;

wire [7:0] recv_tcp_data_cdc_data_out;
cdc_syncfifo #(.DSIZE(8), .ASIZE(3)) cdc_syncfifo_recv_tcp_data
(
    .rdata(recv_tcp_data_cdc_data_out),
    .wfull(recv_tcp_data_wfull),
    .rempty(recv_tcp_data_cdc_fifo_empty),
    .wdata(TCP_RX_DATA),
    .winc(recv_tcp_data_cdc_fifo_write), .wclk(BUS_CLK), .wrst(RESET),
    .rinc(!recv_tcp_data_fifo_full), .rclk(BUS_CLK), .rrst(RESET)
);

always @ (posedge BUS_CLK)
    if(RESET) begin
        TCP_RCV_WRITE_CNT <= 0;
        //TCP_RX_WC <= 0;
    end else if(recv_tcp_data_cdc_fifo_write) begin
        TCP_RCV_WRITE_CNT <= TCP_RCV_WRITE_CNT + 1;
        //TCP_RX_WC <= TCP_RX_WC + 1;
    end else begin
        TCP_RCV_WRITE_CNT <= TCP_RCV_WRITE_CNT;
        //TCP_RX_WC <= 0;
    end

wire RECV_TCP_DATA_FIFO_READ, RECV_TCP_DATA_FIFO_EMPTY;
wire [31:0] RECV_TCP_FIFO_DATA;
fifo_8_to_32 #(.DEPTH(1024)) fifo_recv_tcp_data_i (
    .RST(RESET),
    .CLK(BUS_CLK),
    .WRITE(!recv_tcp_data_cdc_fifo_empty),
    .READ(RECV_TCP_DATA_FIFO_READ),
    .DATA_IN(recv_tcp_data_cdc_data_out),
    .FULL(recv_tcp_data_fifo_full),
    .EMPTY(RECV_TCP_DATA_FIFO_EMPTY),
    .DATA_OUT(RECV_TCP_FIFO_DATA)
);


always @(posedge BUS_CLK)
begin
    if (RESET)
        UDP_WRITE_CNT <= 0;
    else if (BUS_WR && (BUS_ADD >= 2 && BUS_ADD <= 9))
        UDP_WRITE_CNT <= UDP_WRITE_CNT + 1;
    else
        UDP_WRITE_CNT <= UDP_WRITE_CNT;
end

reg [15:0] TCP_WRITE_DLY_CNT;
always @ (posedge BUS_CLK)
    if ((TCP_WRITE_DLY == 0) | RESET)
        TCP_WRITE_DLY_CNT <= 0;
    else if (TCP_WRITE_DLY_CNT == TCP_WRITE_DLY)
        TCP_WRITE_DLY_CNT <= 1;
    else
        TCP_WRITE_DLY_CNT <= TCP_WRITE_DLY_CNT + 1;

reg [31:0] GEN_TCP_DATA;
reg GEN_TCP_DATA_WRITE, GEN_TCP_DATA_WRITE_FF;
always @ (posedge BUS_CLK)
    GEN_TCP_DATA_WRITE_FF <= GEN_TCP_DATA_WRITE;

always @ (posedge BUS_CLK)
    if (TCP_WRITE_DLY == 0 || RESET)
        GEN_TCP_DATA <= 0;
    else if (GEN_TCP_DATA_WRITE_FF)
        GEN_TCP_DATA <= GEN_TCP_DATA + 1;
    else
        GEN_TCP_DATA <= GEN_TCP_DATA;

wire GEN_TCP_DATA_FULL;
wire GEN_TCP_DATA_READ_GRANT;
always @ (posedge BUS_CLK)
    if (RESET)
    begin
        GEN_TCP_DATA_WRITE <= 1'b0;
        TCP_WRITE_CNT <= 0;
        TCP_FAILED_WRITE_CNT <= 0;
    end
    else if (TCP_WRITE_DLY == 0)
    begin
        GEN_TCP_DATA_WRITE <= 1'b0;
        TCP_WRITE_CNT <= TCP_WRITE_CNT;
        TCP_FAILED_WRITE_CNT <= TCP_FAILED_WRITE_CNT;
    end
    else if (TCP_WRITE_DLY == TCP_WRITE_DLY_CNT && !GEN_TCP_DATA_FULL)
    begin
        GEN_TCP_DATA_WRITE <= 1'b1;
        TCP_WRITE_CNT <= TCP_WRITE_CNT + 1;
        TCP_FAILED_WRITE_CNT <= TCP_FAILED_WRITE_CNT;
    end
    else if (TCP_WRITE_DLY == TCP_WRITE_DLY_CNT && GEN_TCP_DATA_FULL)
    begin
        GEN_TCP_DATA_WRITE <= 1'b0;
        TCP_WRITE_CNT <= TCP_WRITE_CNT;
        TCP_FAILED_WRITE_CNT <= TCP_FAILED_WRITE_CNT + 1;
    end
    else
    begin
        GEN_TCP_DATA_WRITE <= 1'b0;
        TCP_WRITE_CNT <= TCP_WRITE_CNT;
        TCP_FAILED_WRITE_CNT <= TCP_FAILED_WRITE_CNT;
    end

wire gen_tcp_data_wfull;
assign GEN_TCP_DATA_FULL = gen_tcp_data_wfull;
wire gen_tcp_data_cdc_fifo_write;
assign gen_tcp_data_cdc_fifo_write = GEN_TCP_DATA_WRITE;
wire gen_tcp_data_fifo_full, gen_tcp_data_cdc_fifo_empty;

wire [31:0] gen_tcp_data_cdc_data_out;
cdc_syncfifo #(.DSIZE(32), .ASIZE(3)) cdc_syncfifo_send_tcp_data_i
(
    .rdata(gen_tcp_data_cdc_data_out),
    .wfull(gen_tcp_data_wfull),
    .rempty(gen_tcp_data_cdc_fifo_empty),
    .wdata(GEN_TCP_DATA),
    .winc(gen_tcp_data_cdc_fifo_write), .wclk(BUS_CLK), .wrst(RESET),
    .rinc(!gen_tcp_data_fifo_full), .rclk(BUS_CLK), .rrst(RESET)
);

wire GEN_TCP_DATA_FIFO_READ, GEN_TCP_DATA_FIFO_EMPTY;
wire [31:0] GEN_TCP_FIFO_DATA;
gerneric_fifo #(
    .DATA_SIZE(32),
    .DEPTH(8)
) fifo_send_tcp_data_i (
    .reset(RESET),
    .clk(BUS_CLK),
    .write(!gen_tcp_data_cdc_fifo_empty),
    .read(GEN_TCP_DATA_FIFO_READ),
    .data_in(gen_tcp_data_cdc_data_out),
    .full(gen_tcp_data_fifo_full),
    .empty(GEN_TCP_DATA_FIFO_EMPTY),
    .data_out(GEN_TCP_FIFO_DATA),
    .size()
);

wire ARB_READY_OUT, ARB_WRITE_OUT;
wire [31:0] ARB_DATA_OUT;
wire [1:0] READ_GRANT;

rrp_arbiter #(
    .WIDTH(2)
) i_rrp_arbiter (
    .RST(RESET),
    .CLK(BUS_CLK),

    .WRITE_REQ({~RECV_TCP_DATA_FIFO_EMPTY, ~GEN_TCP_DATA_FIFO_EMPTY}),
    .HOLD_REQ({2'b0}),
    .DATA_IN({RECV_TCP_FIFO_DATA, GEN_TCP_FIFO_DATA}),
    .READ_GRANT(READ_GRANT),

    .READY_OUT(ARB_READY_OUT),
    .WRITE_OUT(ARB_WRITE_OUT),
    .DATA_OUT(ARB_DATA_OUT)
);

assign GEN_TCP_DATA_FIFO_READ = READ_GRANT[0];
assign RECV_TCP_DATA_FIFO_READ = READ_GRANT[1];
//assign ARB_WRITE_OUT =  GEN_TCP_DATA_WRITE;
//assign ARB_DATA_OUT = GEN_TCP_DATA;

//cdc_fifo is for timing reasons
wire FIFO_FULL;
wire [31:0] cdc_data_out;
wire full_32to8, cdc_fifo_empty;
cdc_syncfifo #(.DSIZE(32), .ASIZE(3)) cdc_syncfifo_i
(
    .rdata(cdc_data_out),
    .wfull(FIFO_FULL),
    .rempty(cdc_fifo_empty),
    .wdata(ARB_DATA_OUT),
    .winc(ARB_WRITE_OUT), .wclk(BUS_CLK), .wrst(RESET),
    .rinc(!full_32to8), .rclk(BUS_CLK), .rrst(RESET)
);
assign ARB_READY_OUT = !FIFO_FULL;

wire FIFO_EMPTY;
fifo_32_to_8 #(.DEPTH(256*1024)) i_data_fifo (
    .RST(RESET),
    .CLK(BUS_CLK),

    .WRITE(!cdc_fifo_empty),
    .READ(TCP_TX_WR),
    .DATA_IN(cdc_data_out),
    .FULL(full_32to8),
    .EMPTY(FIFO_EMPTY),
    .DATA_OUT(TCP_TX_DATA)
);

assign TCP_TX_WR = !TCP_TX_FULL && !FIFO_EMPTY;

wire CLK_1HZ, CE_1HZ;
clock_divider #(
    .DIVISOR(133333333)
) i_clock_divisor_133MHz_to_1Hz (
    .CLK(BUS_CLK),
    .RESET(1'b0),
    .CE(CE_1HZ),
    .CLOCK(CLK_1HZ)
);

wire CLK_3HZ, CE_3HZ;
clock_divider #(
    .DIVISOR(44444444)
) i_clock_divisor_133MHz_to_3Hz (
    .CLK(CLK40),
    .RESET(1'b0),
    .CE(CE_3HZ),
    .CLOCK(CLK_3HZ)
);

wire FIFO_FULL_SYNC;
three_stage_synchronizer #(
    .WIDTH(1)
) three_stage_fifo_full_synchronizer (
    .CLK(BUS_CLK),
    .IN(FIFO_FULL),
    .OUT(FIFO_FULL_SYNC)
);

reg FIFO_WAS_FULL;
always @ (posedge BUS_CLK or posedge FIFO_FULL_SYNC) begin
    if (CE_3HZ || FIFO_FULL_SYNC) begin
        if (FIFO_FULL_SYNC)
            FIFO_WAS_FULL <= 1'b1;
        else
            FIFO_WAS_FULL <= 1'b0;
    end
end

reg FIFO_WAS_ALMOST_EMPTY;
always @ (posedge BUS_CLK or negedge FIFO_FULL_SYNC) begin
    if (CE_3HZ || !FIFO_FULL_SYNC) begin
        if (!FIFO_FULL_SYNC)
            FIFO_WAS_ALMOST_EMPTY <= 1'b1;
        else
            FIFO_WAS_ALMOST_EMPTY <= 1'b0;
    end
end

reg FIFO_FULL_SLOW;
always @ (posedge BUS_CLK or posedge FIFO_WAS_FULL or negedge FIFO_WAS_ALMOST_EMPTY) begin
    if (CE_3HZ || (FIFO_WAS_FULL && !FIFO_WAS_ALMOST_EMPTY)) begin
        if (FIFO_WAS_FULL && !FIFO_WAS_ALMOST_EMPTY)
            FIFO_FULL_SLOW <= 1'b1;
        else if (FIFO_WAS_FULL && !FIFO_FULL_SLOW)
            FIFO_FULL_SLOW <= 1'b1;
        else
            FIFO_FULL_SLOW <= 1'b0;
    end
end

assign LED[7:4] = ~{clock_speed, duplex_status, (|clock_speed & link_status & (GMII_1000M ? CLK_1HZ : CLK_3HZ)) | INVALID};
assign LED[0] = ~CLK_1HZ;
assign LED[1] = ~FIFO_FULL_SLOW;
assign LED[2] = 1'b1;
assign LED[3] = 1'b1;

endmodule
